c1df59abc8abe824c0fd8fd1ec3e3f ����   2 �  weibo4j/org/json/CDL  java/lang/Object <init> ()V Code
  	   LineNumberTable LocalVariableTable this Lweibo4j/org/json/CDL; getValue 2(Lweibo4j/org/json/JSONTokener;)Ljava/lang/String; 
Exceptions  weibo4j/org/json/JSONException
    weibo4j/org/json/JSONTokener   next ()C
     
nextString (C)Ljava/lang/String;
     back !  
  # $  nextTo x Lweibo4j/org/json/JSONTokener; c C StackMapTable rowToJSONArray <(Lweibo4j/org/json/JSONTokener;)Lweibo4j/org/json/JSONArray; - weibo4j/org/json/JSONArray
 , 	
  0  
 , 2 3 4 length ()I
 6 2 7 java/lang/String
 , 9 : ; put 0(Ljava/lang/Object;)Lweibo4j/org/json/JSONArray; = java/lang/StringBuilder ? Bad character '
 < A  B (Ljava/lang/String;)V
 < D E F append (C)Ljava/lang/StringBuilder; H ' (
 < J E K -(Ljava/lang/String;)Ljava/lang/StringBuilder;
 < M E N (I)Ljava/lang/StringBuilder; P ).
 < R S T toString ()Ljava/lang/String;
  V W X syntaxError 4(Ljava/lang/String;)Lweibo4j/org/json/JSONException; ja Lweibo4j/org/json/JSONArray; value Ljava/lang/String; rowToJSONObject Y(Lweibo4j/org/json/JSONArray;Lweibo4j/org/json/JSONTokener;)Lweibo4j/org/json/JSONObject;
  ` * +
 , b c d toJSONObject ;(Lweibo4j/org/json/JSONArray;)Lweibo4j/org/json/JSONObject; names g weibo4j/org/json/JSONObject toJSONArray 0(Ljava/lang/String;)Lweibo4j/org/json/JSONArray;
  A
  l h + string
  o h p X(Lweibo4j/org/json/JSONArray;Lweibo4j/org/json/JSONTokener;)Lweibo4j/org/json/JSONArray; L(Lweibo4j/org/json/JSONArray;Ljava/lang/String;)Lweibo4j/org/json/JSONArray;
  s ] ^ jo Lweibo4j/org/json/JSONObject; rowToString 0(Lweibo4j/org/json/JSONArray;)Ljava/lang/String; y java/lang/StringBuffer
 x 	
 x | E } (C)Ljava/lang/StringBuffer;
 ,  � � opt (I)Ljava/lang/Object;
  R
 6 � � � indexOf (I)I
 x � E � ,(Ljava/lang/String;)Ljava/lang/StringBuffer;
 x R sb Ljava/lang/StringBuffer; i I o Ljava/lang/Object; s
 , � � � optJSONObject  (I)Lweibo4j/org/json/JSONObject;
 f � e � ()Lweibo4j/org/json/JSONArray;
  � v w
 6 � � � valueOf &(Ljava/lang/Object;)Ljava/lang/String;
  � S � L(Lweibo4j/org/json/JSONArray;Lweibo4j/org/json/JSONArray;)Ljava/lang/String;
 f � h � :(Lweibo4j/org/json/JSONArray;)Lweibo4j/org/json/JSONArray; 
SourceFile CDL.java !               /     *� �    
       .             
             �     V*� < ���	����    9          *   "   ,   '   ,   ,   2�*� �*�  �*� *,� "�    
   & 	   :  ;  < < > > A D C H D K F O G        V % &    Q ' (  )   
  � ; 	 * +               p� ,Y� .L*� /M,� +� 1� ,� 5� �+,� 8W*� >,� ��� ���
� � � +�*� <Y>� @� CG� I� LO� I� Q� U�    
   :    R  T  U  V ! X ' Z , [ 2 \ 5 ^ ; _ K ` M b ` c l b    *    p % &    h Y Z   c [ \  , D ' (  )    �  ,�  6�  	 ] ^           g     +� _M,� ,*� a� �    
   
    u  v          e Z      % &    Y Z  )    �  ,@ f 	 h i           6     � Y*� j� k�    
       �         m \   	 h +           3     	*� _*� n�    
       �        	 % &   	 h q           A     *� Y+� j� n�    
       �         e Z      m \  	 h p           �     6*� 
*� 1� �� ,Y� .M*+� rN-� � ,-� 8W���,� 1� �,�    
   .    �  �  �  �  �  � " � ( � + � 2 � 4 �    *    6 e Z     6 % &   ! Y Z    t u  )    �  ,�  f�  	 v w    C     �� xY� zL=� l� 
+,� {W*� ~N-� T-� �:,� �� ="� �� +'� {W+� �W+'� {W� "+"� {W+� �W+"� {W� 
+� �W�*� 1���+
� {W+� ��    
   N    �  �  �  �  �  � " � ( � 2 � < � C � J � T � [ � b � l � s � ~ � � �    4    � Y Z    � � �  
 t � �   U � �  ( K � \  )    �  x
� ;  6�  	 S w           �     /*� �L+� &+� �M,� � <Y,� �� �� @,*� �� I� Q��    
       �  � 
 �  �  � - �         / Y Z    ) t u    e Z  )    � - f 	 S �           �     D*� 
*� 1� �� xY� zM>�  +� �:� ,*� �� �� �W�+� 1���,� ��    
   & 	   �  �  �  �  � ! � &  4 � ?    4    D e Z     D Y Z   / � �   ( � �  !  t u  )    �  x  �    �